`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/10/2022 11:55:32 AM
// Design Name: 
// Module Name: encoder
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module encoder(
    input clk,
    input wire [1023:0] op,
    output reg [9:0] en_op
    );
    
    always @(posedge clk)
      begin
        if (op[1023]==1) en_op = 10'b1111111111;
        else if (op[1021]==1) en_op = 10'b1111111101;
        else if (op[1019]==1) en_op = 10'b1111111011;
        else if (op[1017]==1) en_op = 10'b1111111001;
        else if (op[1015]==1) en_op = 10'b1111110111;
        else if (op[1013]==1) en_op = 10'b1111110101;
        else if (op[1011]==1) en_op = 10'b1111110011;
        else if (op[1009]==1) en_op = 10'b1111110001;
        else if (op[1007]==1) en_op = 10'b1111101111;
        else if (op[1005]==1) en_op = 10'b1111101101;
        else if (op[1003]==1) en_op = 10'b1111101011;
        else if (op[1001]==1) en_op = 10'b1111101001;
        else if (op[999]==1) en_op = 10'b1111100111;
        else if (op[997]==1) en_op = 10'b1111100101;
        else if (op[995]==1) en_op = 10'b1111100011;
        else if (op[993]==1) en_op = 10'b1111100001;
        else if (op[991]==1) en_op = 10'b1111011111;
        else if (op[989]==1) en_op = 10'b1111011101;
        else if (op[987]==1) en_op = 10'b1111011011;
        else if (op[985]==1) en_op = 10'b1111011001;
        else if (op[983]==1) en_op = 10'b1111010111;
        else if (op[981]==1) en_op = 10'b1111010101;
        else if (op[979]==1) en_op = 10'b1111010011;
        else if (op[977]==1) en_op = 10'b1111010001;
        else if (op[975]==1) en_op = 10'b1111001111;
        else if (op[973]==1) en_op = 10'b1111001101;
        else if (op[971]==1) en_op = 10'b1111001011;
        else if (op[969]==1) en_op = 10'b1111001001;
        else if (op[967]==1) en_op = 10'b1111000111;
        else if (op[965]==1) en_op = 10'b1111000101;
        else if (op[963]==1) en_op = 10'b1111000011;
        else if (op[961]==1) en_op = 10'b1111000001;
        else if (op[959]==1) en_op = 10'b1110111111;
        else if (op[957]==1) en_op = 10'b1110111101;
        else if (op[955]==1) en_op = 10'b1110111011;
        else if (op[953]==1) en_op = 10'b1110111001;
        else if (op[951]==1) en_op = 10'b1110110111;
        else if (op[949]==1) en_op = 10'b1110110101;
        else if (op[947]==1) en_op = 10'b1110110011;
        else if (op[945]==1) en_op = 10'b1110110001;
        else if (op[943]==1) en_op = 10'b1110101111;
        else if (op[941]==1) en_op = 10'b1110101101;
        else if (op[939]==1) en_op = 10'b1110101011;
        else if (op[937]==1) en_op = 10'b1110101001;
        else if (op[935]==1) en_op = 10'b1110100111;
        else if (op[933]==1) en_op = 10'b1110100101;
        else if (op[931]==1) en_op = 10'b1110100011;
        else if (op[929]==1) en_op = 10'b1110100001;
        else if (op[927]==1) en_op = 10'b1110011111;
        else if (op[925]==1) en_op = 10'b1110011101;
        else if (op[923]==1) en_op = 10'b1110011011;
        else if (op[921]==1) en_op = 10'b1110011001;
        else if (op[919]==1) en_op = 10'b1110010111;
        else if (op[917]==1) en_op = 10'b1110010101;
        else if (op[915]==1) en_op = 10'b1110010011;
        else if (op[913]==1) en_op = 10'b1110010001;
        else if (op[911]==1) en_op = 10'b1110001111;
        else if (op[909]==1) en_op = 10'b1110001101;
        else if (op[907]==1) en_op = 10'b1110001011;
        else if (op[905]==1) en_op = 10'b1110001001;
        else if (op[903]==1) en_op = 10'b1110000111;
        else if (op[901]==1) en_op = 10'b1110000101;
        else if (op[899]==1) en_op = 10'b1110000011;
        else if (op[897]==1) en_op = 10'b1110000001;
        else if (op[895]==1) en_op = 10'b1101111111;
        else if (op[893]==1) en_op = 10'b1101111101;
        else if (op[891]==1) en_op = 10'b1101111011;
        else if (op[889]==1) en_op = 10'b1101111001;
        else if (op[887]==1) en_op = 10'b1101110111;
        else if (op[885]==1) en_op = 10'b1101110101;
        else if (op[883]==1) en_op = 10'b1101110011;
        else if (op[881]==1) en_op = 10'b1101110001;
        else if (op[879]==1) en_op = 10'b1101101111;
        else if (op[877]==1) en_op = 10'b1101101101;
        else if (op[875]==1) en_op = 10'b1101101011;
        else if (op[873]==1) en_op = 10'b1101101001;
        else if (op[871]==1) en_op = 10'b1101100111;
        else if (op[869]==1) en_op = 10'b1101100101;
        else if (op[867]==1) en_op = 10'b1101100011;
        else if (op[865]==1) en_op = 10'b1101100001;
        else if (op[863]==1) en_op = 10'b1101011111;
        else if (op[861]==1) en_op = 10'b1101011101;
        else if (op[859]==1) en_op = 10'b1101011011;
        else if (op[857]==1) en_op = 10'b1101011001;
        else if (op[855]==1) en_op = 10'b1101010111;
        else if (op[853]==1) en_op = 10'b1101010101;
        else if (op[851]==1) en_op = 10'b1101010011;
        else if (op[849]==1) en_op = 10'b1101010001;
        else if (op[847]==1) en_op = 10'b1101001111;
        else if (op[845]==1) en_op = 10'b1101001101;
        else if (op[843]==1) en_op = 10'b1101001011;
        else if (op[841]==1) en_op = 10'b1101001001;
        else if (op[839]==1) en_op = 10'b1101000111;
        else if (op[837]==1) en_op = 10'b1101000101;
        else if (op[835]==1) en_op = 10'b1101000011;
        else if (op[833]==1) en_op = 10'b1101000001;
        else if (op[831]==1) en_op = 10'b1100111111;
        else if (op[829]==1) en_op = 10'b1100111101;
        else if (op[827]==1) en_op = 10'b1100111011;
        else if (op[825]==1) en_op = 10'b1100111001;
        else if (op[823]==1) en_op = 10'b1100110111;
        else if (op[821]==1) en_op = 10'b1100110101;
        else if (op[819]==1) en_op = 10'b1100110011;
        else if (op[817]==1) en_op = 10'b1100110001;
        else if (op[815]==1) en_op = 10'b1100101111;
        else if (op[813]==1) en_op = 10'b1100101101;
        else if (op[811]==1) en_op = 10'b1100101011;
        else if (op[809]==1) en_op = 10'b1100101001;
        else if (op[807]==1) en_op = 10'b1100100111;
        else if (op[805]==1) en_op = 10'b1100100101;
        else if (op[803]==1) en_op = 10'b1100100011;
        else if (op[801]==1) en_op = 10'b1100100001;
        else if (op[799]==1) en_op = 10'b1100011111;
        else if (op[797]==1) en_op = 10'b1100011101;
        else if (op[795]==1) en_op = 10'b1100011011;
        else if (op[793]==1) en_op = 10'b1100011001;
        else if (op[791]==1) en_op = 10'b1100010111;
        else if (op[789]==1) en_op = 10'b1100010101;
        else if (op[787]==1) en_op = 10'b1100010011;
        else if (op[785]==1) en_op = 10'b1100010001;
        else if (op[783]==1) en_op = 10'b1100001111;
        else if (op[781]==1) en_op = 10'b1100001101;
        else if (op[779]==1) en_op = 10'b1100001011;
        else if (op[777]==1) en_op = 10'b1100001001;
        else if (op[775]==1) en_op = 10'b1100000111;
        else if (op[773]==1) en_op = 10'b1100000101;
        else if (op[771]==1) en_op = 10'b1100000011;
        else if (op[769]==1) en_op = 10'b1100000001;
        else if (op[767]==1) en_op = 10'b1011111111;
        else if (op[765]==1) en_op = 10'b1011111101;
        else if (op[763]==1) en_op = 10'b1011111011;
        else if (op[761]==1) en_op = 10'b1011111001;
        else if (op[759]==1) en_op = 10'b1011110111;
        else if (op[757]==1) en_op = 10'b1011110101;
        else if (op[755]==1) en_op = 10'b1011110011;
        else if (op[753]==1) en_op = 10'b1011110001;
        else if (op[751]==1) en_op = 10'b1011101111;
        else if (op[749]==1) en_op = 10'b1011101101;
        else if (op[747]==1) en_op = 10'b1011101011;
        else if (op[745]==1) en_op = 10'b1011101001;
        else if (op[743]==1) en_op = 10'b1011100111;
        else if (op[741]==1) en_op = 10'b1011100101;
        else if (op[739]==1) en_op = 10'b1011100011;
        else if (op[737]==1) en_op = 10'b1011100001;
        else if (op[735]==1) en_op = 10'b1011011111;
        else if (op[733]==1) en_op = 10'b1011011101;
        else if (op[731]==1) en_op = 10'b1011011011;
        else if (op[729]==1) en_op = 10'b1011011001;
        else if (op[727]==1) en_op = 10'b1011010111;
        else if (op[725]==1) en_op = 10'b1011010101;
        else if (op[723]==1) en_op = 10'b1011010011;
        else if (op[721]==1) en_op = 10'b1011010001;
        else if (op[719]==1) en_op = 10'b1011001111;
        else if (op[717]==1) en_op = 10'b1011001101;
        else if (op[715]==1) en_op = 10'b1011001011;
        else if (op[713]==1) en_op = 10'b1011001001;
        else if (op[711]==1) en_op = 10'b1011000111;
        else if (op[709]==1) en_op = 10'b1011000101;
        else if (op[707]==1) en_op = 10'b1011000011;
        else if (op[705]==1) en_op = 10'b1011000001;
        else if (op[703]==1) en_op = 10'b1010111111;
        else if (op[701]==1) en_op = 10'b1010111101;
        else if (op[699]==1) en_op = 10'b1010111011;
        else if (op[697]==1) en_op = 10'b1010111001;
        else if (op[695]==1) en_op = 10'b1010110111;
        else if (op[693]==1) en_op = 10'b1010110101;
        else if (op[691]==1) en_op = 10'b1010110011;
        else if (op[689]==1) en_op = 10'b1010110001;
        else if (op[687]==1) en_op = 10'b1010101111;
        else if (op[685]==1) en_op = 10'b1010101101;
        else if (op[683]==1) en_op = 10'b1010101011;
        else if (op[681]==1) en_op = 10'b1010101001;
        else if (op[679]==1) en_op = 10'b1010100111;
        else if (op[677]==1) en_op = 10'b1010100101;
        else if (op[675]==1) en_op = 10'b1010100011;
        else if (op[673]==1) en_op = 10'b1010100001;
        else if (op[671]==1) en_op = 10'b1010011111;
        else if (op[669]==1) en_op = 10'b1010011101;
        else if (op[667]==1) en_op = 10'b1010011011;
        else if (op[665]==1) en_op = 10'b1010011001;
        else if (op[663]==1) en_op = 10'b1010010111;
        else if (op[661]==1) en_op = 10'b1010010101;
        else if (op[659]==1) en_op = 10'b1010010011;
        else if (op[657]==1) en_op = 10'b1010010001;
        else if (op[655]==1) en_op = 10'b1010001111;
        else if (op[653]==1) en_op = 10'b1010001101;
        else if (op[651]==1) en_op = 10'b1010001011;
        else if (op[649]==1) en_op = 10'b1010001001;
        else if (op[647]==1) en_op = 10'b1010000111;
        else if (op[645]==1) en_op = 10'b1010000101;
        else if (op[643]==1) en_op = 10'b1010000011;
        else if (op[641]==1) en_op = 10'b1010000001;
        else if (op[639]==1) en_op = 10'b1001111111;
        else if (op[637]==1) en_op = 10'b1001111101;
        else if (op[635]==1) en_op = 10'b1001111011;
        else if (op[633]==1) en_op = 10'b1001111001;
        else if (op[631]==1) en_op = 10'b1001110111;
        else if (op[629]==1) en_op = 10'b1001110101;
        else if (op[627]==1) en_op = 10'b1001110011;
        else if (op[625]==1) en_op = 10'b1001110001;
        else if (op[623]==1) en_op = 10'b1001101111;
        else if (op[621]==1) en_op = 10'b1001101101;
        else if (op[619]==1) en_op = 10'b1001101011;
        else if (op[617]==1) en_op = 10'b1001101001;
        else if (op[615]==1) en_op = 10'b1001100111;
        else if (op[613]==1) en_op = 10'b1001100101;
        else if (op[611]==1) en_op = 10'b1001100011;
        else if (op[609]==1) en_op = 10'b1001100001;
        else if (op[607]==1) en_op = 10'b1001011111;
        else if (op[605]==1) en_op = 10'b1001011101;
        else if (op[603]==1) en_op = 10'b1001011011;
        else if (op[601]==1) en_op = 10'b1001011001;
        else if (op[599]==1) en_op = 10'b1001010111;
        else if (op[597]==1) en_op = 10'b1001010101;
        else if (op[595]==1) en_op = 10'b1001010011;
        else if (op[593]==1) en_op = 10'b1001010001;
        else if (op[591]==1) en_op = 10'b1001001111;
        else if (op[589]==1) en_op = 10'b1001001101;
        else if (op[587]==1) en_op = 10'b1001001011;
        else if (op[585]==1) en_op = 10'b1001001001;
        else if (op[583]==1) en_op = 10'b1001000111;
        else if (op[581]==1) en_op = 10'b1001000101;
        else if (op[579]==1) en_op = 10'b1001000011;
        else if (op[577]==1) en_op = 10'b1001000001;
        else if (op[575]==1) en_op = 10'b1000111111;
        else if (op[573]==1) en_op = 10'b1000111101;
        else if (op[571]==1) en_op = 10'b1000111011;
        else if (op[569]==1) en_op = 10'b1000111001;
        else if (op[567]==1) en_op = 10'b1000110111;
        else if (op[565]==1) en_op = 10'b1000110101;
        else if (op[563]==1) en_op = 10'b1000110011;
        else if (op[561]==1) en_op = 10'b1000110001;
        else if (op[559]==1) en_op = 10'b1000101111;
        else if (op[557]==1) en_op = 10'b1000101101;
        else if (op[555]==1) en_op = 10'b1000101011;
        else if (op[553]==1) en_op = 10'b1000101001;
        else if (op[551]==1) en_op = 10'b1000100111;
        else if (op[549]==1) en_op = 10'b1000100101;
        else if (op[547]==1) en_op = 10'b1000100011;
        else if (op[545]==1) en_op = 10'b1000100001;
        else if (op[543]==1) en_op = 10'b1000011111;
        else if (op[541]==1) en_op = 10'b1000011101;
        else if (op[539]==1) en_op = 10'b1000011011;
        else if (op[537]==1) en_op = 10'b1000011001;
        else if (op[535]==1) en_op = 10'b1000010111;
        else if (op[533]==1) en_op = 10'b1000010101;
        else if (op[531]==1) en_op = 10'b1000010011;
        else if (op[529]==1) en_op = 10'b1000010001;
        else if (op[527]==1) en_op = 10'b1000001111;
        else if (op[525]==1) en_op = 10'b1000001101;
        else if (op[523]==1) en_op = 10'b1000001011;
        else if (op[521]==1) en_op = 10'b1000001001;
        else if (op[519]==1) en_op = 10'b1000000111;
        else if (op[517]==1) en_op = 10'b1000000101;
        else if (op[515]==1) en_op = 10'b1000000011;
        else if (op[513]==1) en_op = 10'b1000000001;
        else if (op[511]==1) en_op = 10'b0111111111;
        else if (op[509]==1) en_op = 10'b0111111101;
        else if (op[507]==1) en_op = 10'b0111111011;
        else if (op[505]==1) en_op = 10'b0111111001;
        else if (op[503]==1) en_op = 10'b0111110111;
        else if (op[501]==1) en_op = 10'b0111110101;
        else if (op[499]==1) en_op = 10'b0111110011;
        else if (op[497]==1) en_op = 10'b0111110001;
        else if (op[495]==1) en_op = 10'b0111101111;
        else if (op[493]==1) en_op = 10'b0111101101;
        else if (op[491]==1) en_op = 10'b0111101011;
        else if (op[489]==1) en_op = 10'b0111101001;
        else if (op[487]==1) en_op = 10'b0111100111;
        else if (op[485]==1) en_op = 10'b0111100101;
        else if (op[483]==1) en_op = 10'b0111100011;
        else if (op[481]==1) en_op = 10'b0111100001;
        else if (op[479]==1) en_op = 10'b0111011111;
        else if (op[477]==1) en_op = 10'b0111011101;
        else if (op[475]==1) en_op = 10'b0111011011;
        else if (op[473]==1) en_op = 10'b0111011001;
        else if (op[471]==1) en_op = 10'b0111010111;
        else if (op[469]==1) en_op = 10'b0111010101;
        else if (op[467]==1) en_op = 10'b0111010011;
        else if (op[465]==1) en_op = 10'b0111010001;
        else if (op[463]==1) en_op = 10'b0111001111;
        else if (op[461]==1) en_op = 10'b0111001101;
        else if (op[459]==1) en_op = 10'b0111001011;
        else if (op[457]==1) en_op = 10'b0111001001;
        else if (op[455]==1) en_op = 10'b0111000111;
        else if (op[453]==1) en_op = 10'b0111000101;
        else if (op[451]==1) en_op = 10'b0111000011;
        else if (op[449]==1) en_op = 10'b0111000001;
        else if (op[447]==1) en_op = 10'b0110111111;
        else if (op[445]==1) en_op = 10'b0110111101;
        else if (op[443]==1) en_op = 10'b0110111011;
        else if (op[441]==1) en_op = 10'b0110111001;
        else if (op[439]==1) en_op = 10'b0110110111;
        else if (op[437]==1) en_op = 10'b0110110101;
        else if (op[435]==1) en_op = 10'b0110110011;
        else if (op[433]==1) en_op = 10'b0110110001;
        else if (op[431]==1) en_op = 10'b0110101111;
        else if (op[429]==1) en_op = 10'b0110101101;
        else if (op[427]==1) en_op = 10'b0110101011;
        else if (op[425]==1) en_op = 10'b0110101001;
        else if (op[423]==1) en_op = 10'b0110100111;
        else if (op[421]==1) en_op = 10'b0110100101;
        else if (op[419]==1) en_op = 10'b0110100011;
        else if (op[417]==1) en_op = 10'b0110100001;
        else if (op[415]==1) en_op = 10'b0110011111;
        else if (op[413]==1) en_op = 10'b0110011101;
        else if (op[411]==1) en_op = 10'b0110011011;
        else if (op[409]==1) en_op = 10'b0110011001;
        else if (op[407]==1) en_op = 10'b0110010111;
        else if (op[405]==1) en_op = 10'b0110010101;
        else if (op[403]==1) en_op = 10'b0110010011;
        else if (op[401]==1) en_op = 10'b0110010001;
        else if (op[399]==1) en_op = 10'b0110001111;
        else if (op[397]==1) en_op = 10'b0110001101;
        else if (op[395]==1) en_op = 10'b0110001011;
        else if (op[393]==1) en_op = 10'b0110001001;
        else if (op[391]==1) en_op = 10'b0110000111;
        else if (op[389]==1) en_op = 10'b0110000101;
        else if (op[387]==1) en_op = 10'b0110000011;
        else if (op[385]==1) en_op = 10'b0110000001;
        else if (op[383]==1) en_op = 10'b0101111111;
        else if (op[381]==1) en_op = 10'b0101111101;
        else if (op[379]==1) en_op = 10'b0101111011;
        else if (op[377]==1) en_op = 10'b0101111001;
        else if (op[375]==1) en_op = 10'b0101110111;
        else if (op[373]==1) en_op = 10'b0101110101;
        else if (op[371]==1) en_op = 10'b0101110011;
        else if (op[369]==1) en_op = 10'b0101110001;
        else if (op[367]==1) en_op = 10'b0101101111;
        else if (op[365]==1) en_op = 10'b0101101101;
        else if (op[363]==1) en_op = 10'b0101101011;
        else if (op[361]==1) en_op = 10'b0101101001;
        else if (op[359]==1) en_op = 10'b0101100111;
        else if (op[357]==1) en_op = 10'b0101100101;
        else if (op[355]==1) en_op = 10'b0101100011;
        else if (op[353]==1) en_op = 10'b0101100001;
        else if (op[351]==1) en_op = 10'b0101011111;
        else if (op[349]==1) en_op = 10'b0101011101;
        else if (op[347]==1) en_op = 10'b0101011011;
        else if (op[345]==1) en_op = 10'b0101011001;
        else if (op[343]==1) en_op = 10'b0101010111;
        else if (op[341]==1) en_op = 10'b0101010101;
        else if (op[339]==1) en_op = 10'b0101010011;
        else if (op[337]==1) en_op = 10'b0101010001;
        else if (op[335]==1) en_op = 10'b0101001111;
        else if (op[333]==1) en_op = 10'b0101001101;
        else if (op[331]==1) en_op = 10'b0101001011;
        else if (op[329]==1) en_op = 10'b0101001001;
        else if (op[327]==1) en_op = 10'b0101000111;
        else if (op[325]==1) en_op = 10'b0101000101;
        else if (op[323]==1) en_op = 10'b0101000011;
        else if (op[321]==1) en_op = 10'b0101000001;
        else if (op[319]==1) en_op = 10'b0100111111;
        else if (op[317]==1) en_op = 10'b0100111101;
        else if (op[315]==1) en_op = 10'b0100111011;
        else if (op[313]==1) en_op = 10'b0100111001;
        else if (op[311]==1) en_op = 10'b0100110111;
        else if (op[309]==1) en_op = 10'b0100110101;
        else if (op[307]==1) en_op = 10'b0100110011;
        else if (op[305]==1) en_op = 10'b0100110001;
        else if (op[303]==1) en_op = 10'b0100101111;
        else if (op[301]==1) en_op = 10'b0100101101;
        else if (op[299]==1) en_op = 10'b0100101011;
        else if (op[297]==1) en_op = 10'b0100101001;
        else if (op[295]==1) en_op = 10'b0100100111;
        else if (op[293]==1) en_op = 10'b0100100101;
        else if (op[291]==1) en_op = 10'b0100100011;
        else if (op[289]==1) en_op = 10'b0100100001;
        else if (op[287]==1) en_op = 10'b0100011111;
        else if (op[285]==1) en_op = 10'b0100011101;
        else if (op[283]==1) en_op = 10'b0100011011;
        else if (op[281]==1) en_op = 10'b0100011001;
        else if (op[279]==1) en_op = 10'b0100010111;
        else if (op[277]==1) en_op = 10'b0100010101;
        else if (op[275]==1) en_op = 10'b0100010011;
        else if (op[273]==1) en_op = 10'b0100010001;
        else if (op[271]==1) en_op = 10'b0100001111;
        else if (op[269]==1) en_op = 10'b0100001101;
        else if (op[267]==1) en_op = 10'b0100001011;
        else if (op[265]==1) en_op = 10'b0100001001;
        else if (op[263]==1) en_op = 10'b0100000111;
        else if (op[261]==1) en_op = 10'b0100000101;
        else if (op[259]==1) en_op = 10'b0100000011;
        else if (op[257]==1) en_op = 10'b0100000001;
        else if (op[255]==1) en_op = 10'b0011111111;
        else if (op[253]==1) en_op = 10'b0011111101;
        else if (op[251]==1) en_op = 10'b0011111011;
        else if (op[249]==1) en_op = 10'b0011111001;
        else if (op[247]==1) en_op = 10'b0011110111;
        else if (op[245]==1) en_op = 10'b0011110101;
        else if (op[243]==1) en_op = 10'b0011110011;
        else if (op[241]==1) en_op = 10'b0011110001;
        else if (op[239]==1) en_op = 10'b0011101111;
        else if (op[237]==1) en_op = 10'b0011101101;
        else if (op[235]==1) en_op = 10'b0011101011;
        else if (op[233]==1) en_op = 10'b0011101001;
        else if (op[231]==1) en_op = 10'b0011100111;
        else if (op[229]==1) en_op = 10'b0011100101;
        else if (op[227]==1) en_op = 10'b0011100011;
        else if (op[225]==1) en_op = 10'b0011100001;
        else if (op[223]==1) en_op = 10'b0011011111;
        else if (op[221]==1) en_op = 10'b0011011101;
        else if (op[219]==1) en_op = 10'b0011011011;
        else if (op[217]==1) en_op = 10'b0011011001;
        else if (op[215]==1) en_op = 10'b0011010111;
        else if (op[213]==1) en_op = 10'b0011010101;
        else if (op[211]==1) en_op = 10'b0011010011;
        else if (op[209]==1) en_op = 10'b0011010001;
        else if (op[207]==1) en_op = 10'b0011001111;
        else if (op[205]==1) en_op = 10'b0011001101;
        else if (op[203]==1) en_op = 10'b0011001011;
        else if (op[201]==1) en_op = 10'b0011001001;
        else if (op[199]==1) en_op = 10'b0011000111;
        else if (op[197]==1) en_op = 10'b0011000101;
        else if (op[195]==1) en_op = 10'b0011000011;
        else if (op[193]==1) en_op = 10'b0011000001;
        else if (op[191]==1) en_op = 10'b0010111111;
        else if (op[189]==1) en_op = 10'b0010111101;
        else if (op[187]==1) en_op = 10'b0010111011;
        else if (op[185]==1) en_op = 10'b0010111001;
        else if (op[183]==1) en_op = 10'b0010110111;
        else if (op[181]==1) en_op = 10'b0010110101;
        else if (op[179]==1) en_op = 10'b0010110011;
        else if (op[177]==1) en_op = 10'b0010110001;
        else if (op[175]==1) en_op = 10'b0010101111;
        else if (op[173]==1) en_op = 10'b0010101101;
        else if (op[171]==1) en_op = 10'b0010101011;
        else if (op[169]==1) en_op = 10'b0010101001;
        else if (op[167]==1) en_op = 10'b0010100111;
        else if (op[165]==1) en_op = 10'b0010100101;
        else if (op[163]==1) en_op = 10'b0010100011;
        else if (op[161]==1) en_op = 10'b0010100001;
        else if (op[159]==1) en_op = 10'b0010011111;
        else if (op[157]==1) en_op = 10'b0010011101;
        else if (op[155]==1) en_op = 10'b0010011011;
        else if (op[153]==1) en_op = 10'b0010011001;
        else if (op[151]==1) en_op = 10'b0010010111;
        else if (op[149]==1) en_op = 10'b0010010101;
        else if (op[147]==1) en_op = 10'b0010010011;
        else if (op[145]==1) en_op = 10'b0010010001;
        else if (op[143]==1) en_op = 10'b0010001111;
        else if (op[141]==1) en_op = 10'b0010001101;
        else if (op[139]==1) en_op = 10'b0010001011;
        else if (op[137]==1) en_op = 10'b0010001001;
        else if (op[135]==1) en_op = 10'b0010000111;
        else if (op[133]==1) en_op = 10'b0010000101;
        else if (op[131]==1) en_op = 10'b0010000011;
        else if (op[129]==1) en_op = 10'b0010000001;
        else if (op[127]==1) en_op = 10'b0001111111;
        else if (op[125]==1) en_op = 10'b0001111101;
        else if (op[123]==1) en_op = 10'b0001111011;
        else if (op[121]==1) en_op = 10'b0001111001;
        else if (op[119]==1) en_op = 10'b0001110111;
        else if (op[117]==1) en_op = 10'b0001110101;
        else if (op[115]==1) en_op = 10'b0001110011;
        else if (op[113]==1) en_op = 10'b0001110001;
        else if (op[111]==1) en_op = 10'b0001101111;
        else if (op[109]==1) en_op = 10'b0001101101;
        else if (op[107]==1) en_op = 10'b0001101011;
        else if (op[105]==1) en_op = 10'b0001101001;
        else if (op[103]==1) en_op = 10'b0001100111;
        else if (op[101]==1) en_op = 10'b0001100101;
        else if (op[99]==1) en_op = 10'b0001100011;
        else if (op[97]==1) en_op = 10'b0001100001;
        else if (op[95]==1) en_op = 10'b0001011111;
        else if (op[93]==1) en_op = 10'b0001011101;
        else if (op[91]==1) en_op = 10'b0001011011;
        else if (op[89]==1) en_op = 10'b0001011001;
        else if (op[87]==1) en_op = 10'b0001010111;
        else if (op[85]==1) en_op = 10'b0001010101;
        else if (op[83]==1) en_op = 10'b0001010011;
        else if (op[81]==1) en_op = 10'b0001010001;
        else if (op[79]==1) en_op = 10'b0001001111;
        else if (op[77]==1) en_op = 10'b0001001101;
        else if (op[75]==1) en_op = 10'b0001001011;
        else if (op[73]==1) en_op = 10'b0001001001;
        else if (op[71]==1) en_op = 10'b0001000111;
        else if (op[69]==1) en_op = 10'b0001000101;
        else if (op[67]==1) en_op = 10'b0001000011;
        else if (op[65]==1) en_op = 10'b0001000001;
        else if (op[63]==1) en_op = 10'b0000111111;
        else if (op[61]==1) en_op = 10'b0000111101;
        else if (op[59]==1) en_op = 10'b0000111011;
        else if (op[57]==1) en_op = 10'b0000111001;
        else if (op[55]==1) en_op = 10'b0000110111;
        else if (op[53]==1) en_op = 10'b0000110101;
        else if (op[51]==1) en_op = 10'b0000110011;
        else if (op[49]==1) en_op = 10'b0000110001;
        else if (op[47]==1) en_op = 10'b0000101111;
        else if (op[45]==1) en_op = 10'b0000101101;
        else if (op[43]==1) en_op = 10'b0000101011;
        else if (op[41]==1) en_op = 10'b0000101001;
        else if (op[39]==1) en_op = 10'b0000100111;
        else if (op[37]==1) en_op = 10'b0000100101;
        else if (op[35]==1) en_op = 10'b0000100011;
        else if (op[33]==1) en_op = 10'b0000100001;
        else if (op[31]==1) en_op = 10'b0000011111;
        else if (op[29]==1) en_op = 10'b0000011101;
        else if (op[27]==1) en_op = 10'b0000011011;
        else if (op[25]==1) en_op = 10'b0000011001;
        else if (op[23]==1) en_op = 10'b0000010111;
        else if (op[21]==1) en_op = 10'b0000010101;
        else if (op[19]==1) en_op = 10'b0000010011;
        else if (op[17]==1) en_op = 10'b0000010001;
        else if (op[15]==1) en_op = 10'b0000001111;
        else if (op[13]==1) en_op = 10'b0000001101;
        else if (op[11]==1) en_op = 10'b0000001011;
        else if (op[9]==1) en_op = 10'b0000001001;
        else if (op[7]==1) en_op = 10'b0000000111;
        else if (op[5]==1) en_op = 10'b0000000101;
        else if (op[3]==1) en_op = 10'b0000000011;
        else if (op[1]==1) en_op = 10'b0000000001;
        else
        en_op = 10'b0000000000;
      end

endmodule
